module maj_vote(
input logic             x0_i,
input logic             x1_i,
input logic             x2_i,
output logic            y_o
);

endmodule
